<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-147.938,39.1654,-56.1383,-6.20957</PageViewport>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>-98.5,63</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>-98.5,59.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>-78,61</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>-101,64.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>-101.5,60</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AE_OR2</type>
<position>-90,61.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>BE_NOR2</type>
<position>-86,53</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>-95,54.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>-95,51.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>-78,53</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND3</type>
<position>-65.5,40.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<input>
<ID>IN_2</ID>16 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>-74,43</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>-73.5,41</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>-73.5,38.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>-53.5,40.5</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>-118,34.5</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>-118,43.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>-118,38.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>-80.5,41.5</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>-103.5,48.5</position>
<gparam>LABEL_TEXT F=x+y'z</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>-122,44.5</position>
<gparam>LABEL_TEXT x</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_AND2</type>
<position>-100,37.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_INVERTER</type>
<position>-110.5,38.5</position>
<input>
<ID>IN_0</ID>22 </input>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>58</ID>
<type>AE_OR2</type>
<position>-91.5,44.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>-120.5,45.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>-121,39.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>-121,35</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>-106,41.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>-129.5,19</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>-129.5,15</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>-130,-2.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>-123.5,18.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>-123.5,14.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_TOGGLE</type>
<position>-125.5,-3.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_AND2</type>
<position>-111.5,18.5</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_AND2</type>
<position>-112,13</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_AND2</type>
<position>-111.5,7.5</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_AND2</type>
<position>-111.5,1</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-94.5,62.5,-94.5,63</points>
<intersection>62.5 1</intersection>
<intersection>63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-94.5,62.5,-93,62.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-94.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-96.5,63,-94.5,63</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-94.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-94.5,59.5,-94.5,60.5</points>
<intersection>59.5 2</intersection>
<intersection>60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-94.5,60.5,-93,60.5</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>-94.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-96.5,59.5,-94.5,59.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-94.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-83,61,-83,61.5</points>
<intersection>61 1</intersection>
<intersection>61.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-83,61,-79,61</points>
<connection>
<GID>12</GID>
<name>N_in0</name></connection>
<intersection>-83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-87,61.5,-83,61.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>-83 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-91,54,-91,54.5</points>
<intersection>54 1</intersection>
<intersection>54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-91,54,-89,54</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-91 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-93,54.5,-91,54.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-91 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-91,51.5,-91,52</points>
<intersection>51.5 2</intersection>
<intersection>52 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-91,52,-89,52</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-91 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-93,51.5,-91,51.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-91 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-83,53,-79,53</points>
<connection>
<GID>28</GID>
<name>N_in0</name></connection>
<connection>
<GID>22</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-72,42.5,-68.5,42.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-72 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-72,42.5,-72,43</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>42.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71.5,40.5,-68.5,40.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>-71.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-71.5,40.5,-71.5,41</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>40.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71.5,38.5,-68.5,38.5</points>
<connection>
<GID>30</GID>
<name>IN_2</name></connection>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-62.5,40.5,-54.5,40.5</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<connection>
<GID>38</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,38.5,-113.5,38.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109.5,34.5,-109.5,36.5</points>
<intersection>34.5 2</intersection>
<intersection>36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-109.5,36.5,-103,36.5</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>-109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116,34.5,-109.5,34.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-107.5,38.5,-103,38.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-105,43.5,-105,45.5</points>
<intersection>43.5 2</intersection>
<intersection>45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-105,45.5,-94.5,45.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-105 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116,43.5,-105,43.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>-105 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-95.5,37.5,-95.5,43.5</points>
<intersection>37.5 2</intersection>
<intersection>43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-95.5,43.5,-94.5,43.5</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>-95.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-97,37.5,-95.5,37.5</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>-95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-85,41.5,-85,44.5</points>
<intersection>41.5 1</intersection>
<intersection>44.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-85,41.5,-81.5,41.5</points>
<connection>
<GID>48</GID>
<name>N_in0</name></connection>
<intersection>-85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-88.5,44.5,-85,44.5</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<intersection>-85 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>